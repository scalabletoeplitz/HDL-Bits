module top_module(
    output zero
);// Module body starts after semicolon

    assign zero = 2'b00;
    
endmodule
